// ****************************************************************************
// ****************************************************************************
// Copyright SoC Design Research Group, All rights reservxd.
// Electronics and Telecommunications Research Institute (ETRI)
// 
// THESE DOCUMENTS CONTAIN CONFIDENTIAL INFORMATION AND KNOWLEDGE
// WHICH IS THE PROPERTY OF ETRI. NO PART OF THIS PUBLICATION IS
// TO BE USED FOR ANY OTHER PURPOSE, AND THESE ARE NOT TO BE
// REPRODUCED, COPIED, DISCLOSED, TRANSMITTED, STORED IN A RETRIEVAL
// SYSTEM OR TRANSLATED INTO ANY OTHER HUMAN OR COMPUTER LANGUAGE,
// IN ANY FORM, BY ANY MEANS, IN WHOLE OR IN PART, WITHOUT THE
// COMPLETE PRIOR WRITTEN PERMISSION OF ETRI.
// ****************************************************************************
// 2025-11-05
// Kyuseung Han (han@etri.re.kr)
// ****************************************************************************
// ****************************************************************************
`ifndef DCA_GDEF_51
`define DCA_GDEF_51

`define DCA_GDEF_24 544
`define DCA_GDEF_46 0

`define DCA_GDEF_16 32
`define DCA_GDEF_01 0

`define DCA_GDEF_13 32
`define DCA_GDEF_32 0

`define DCA_GDEF_15 16
`define DCA_GDEF_21 0
`define DCA_GDEF_48 1
`define DCA_GDEF_18 2
`define DCA_GDEF_19 4
`define DCA_GDEF_35 8
`define DCA_GDEF_25 16
`define DCA_GDEF_60 32
`define DCA_GDEF_49 64
`define DCA_GDEF_29 128
`define DCA_GDEF_30 256
`define DCA_GDEF_52 512
`define DCA_GDEF_28 1024
`define DCA_GDEF_45 2048
`define DCA_GDEF_14 4096
`define DCA_GDEF_47 8192
`define DCA_GDEF_41 16384
`define DCA_GDEF_26 32768
`define DCA_GDEF_39 0
`define DCA_GDEF_02 1
`define DCA_GDEF_10 2
`define DCA_GDEF_40 3
`define DCA_GDEF_31 4
`define DCA_GDEF_00 5
`define DCA_GDEF_54 6
`define DCA_GDEF_36 7
`define DCA_GDEF_22 8
`define DCA_GDEF_06 9
`define DCA_GDEF_50 10
`define DCA_GDEF_27 11
`define DCA_GDEF_55 12
`define DCA_GDEF_43 13
`define DCA_GDEF_58 14
`define DCA_GDEF_42 15
`define DCA_GDEF_05 0

`define DCA_GDEF_44 8
`define DCA_GDEF_20 0

`define DCA_GDEF_33 512
`define DCA_GDEF_23 0

`define DCA_GDEF_12 4
`define DCA_GDEF_53 0

`define DCA_GDEF_17 4
`define DCA_GDEF_04 0

`define DCA_GDEF_11 32
`define DCA_GDEF_38 0

`define DCA_GDEF_34 32
`define DCA_GDEF_08 0

`define DCA_GDEF_37 2
`define DCA_GDEF_56 0
`define DCA_GDEF_07 1
`define DCA_GDEF_59 2
`define DCA_GDEF_57 0
`define DCA_GDEF_09 1
`define DCA_GDEF_03 0

`endif