// ****************************************************************************
// ****************************************************************************
// Copyright SoC Design Research Group, All rights reserved.
// Electronics and Telecommunications Research Institute (ETRI)
// 
// THESE DOCUMENTS CONTAIN CONFIDENTIAL INFORMATION AND KNOWLEDGE
// WHICH IS THE PROPERTY OF ETRI. NO PART OF THIS PUBLICATION IS
// TO BE USED FOR ANY OTHER PURPOSE, AND THESE ARE NOT TO BE
// REPRODUCED, COPIED, DISCLOSED, TRANSMITTED, STORED IN A RETRIEVAL
// SYSTEM OR TRANSLATED INTO ANY OTHER HUMAN OR COMPUTER LANGUAGE,
// IN ANY FORM, BY ANY MEANS, IN WHOLE OR IN PART, WITHOUT THE
// COMPLETE PRIOR WRITTEN PERMISSION OF ETRI.
// ****************************************************************************
// 2025-10-31
// Kyuseung Han (han@etri.re.kr)
// ****************************************************************************
// ****************************************************************************

`include "ervp_platform_controller_memorymap_offset.vh"
`include "ervp_external_peri_group_memorymap_offset.vh"
`include "memorymap_info.vh"
`include "ervp_global.vh"
`include "platform_info.vh"
`include "munoc_network_include.vh"

module FSD_V1
(
	xa_p0,
	xa_n0,
	external_clk_0,
	external_clk_0_pair,
	external_rstnn,
	led_list,
	switch_slide_readymade_0,
	gpio0,
	gpio1,
	gpio2,
	gpio3,
	gpio4,
	pjtag_rtck,
	pjtag_rtrstnn,
	pjtag_rtms,
	pjtag_rtdi,
	pjtag_rtdo,
	printf_tx,
	printf_rx
	`include "slow_dram_cell_port_dec.vh"
);


input wire xa_p0;
input wire xa_n0;
input wire external_clk_0;
input wire external_clk_0_pair;
input wire external_rstnn;
output wire [((1)*(1))-1:0] led_list;
inout wire switch_slide_readymade_0;
inout wire gpio0;
inout wire gpio1;
inout wire gpio2;
inout wire gpio3;
inout wire gpio4;
input wire pjtag_rtck;
input wire pjtag_rtrstnn;
input wire pjtag_rtms;
input wire pjtag_rtdi;
output wire pjtag_rtdo;
output wire printf_tx;
input wire printf_rx;

`include "slow_dram_cell_port_def.vh"


wire clk_system;
wire clk_dca_core;
wire clk_core;
wire clk_system_external;
wire clk_system_debug;
wire clk_local_access;
wire clk_process_000;
wire clk_process_001;
wire clk_dram_if;
wire clk_dram_sys;
wire clk_dram_ref;
wire clk_noc;
wire gclk_system;
wire gclk_dca_core;
wire gclk_core;
wire gclk_system_external;
wire gclk_system_debug;
wire gclk_local_access;
wire gclk_process_000;
wire gclk_process_001;
wire gclk_noc;
wire tick_1us;
wire tick_62d5ms;
wire tick_gpio;
wire spi_common_sclk;
wire spi_common_sdq0;
wire global_rstnn;
wire global_rstpp;
wire [(9)-1:0] rstnn_seqeunce;
wire [(9)-1:0] rstpp_seqeunce;
wire rstnn_user;
wire rstpp_user;
wire i_rtl_clk_system;
wire i_rtl_clk_dca_core;
wire i_rtl_clk_core;
wire i_rtl_clk_system_external;
wire i_rtl_clk_system_debug;
wire i_rtl_clk_local_access;
wire i_rtl_clk_process_000;
wire i_rtl_clk_process_001;
wire i_rtl_clk_dram_if;
wire i_rtl_clk_dram_sys;
wire i_rtl_clk_dram_ref;
wire i_rtl_clk_noc;
wire i_rtl_gclk_system;
wire i_rtl_gclk_dca_core;
wire i_rtl_gclk_core;
wire i_rtl_gclk_system_external;
wire i_rtl_gclk_system_debug;
wire i_rtl_gclk_local_access;
wire i_rtl_gclk_process_000;
wire i_rtl_gclk_process_001;
wire i_rtl_gclk_noc;
wire i_rtl_tick_1us;
wire i_rtl_tick_62d5ms;
wire i_rtl_tick_gpio;
wire i_rtl_spi_common_sclk;
wire i_rtl_spi_common_sdq0;
wire i_rtl_external_rstnn;
wire i_rtl_global_rstnn;
wire i_rtl_global_rstpp;
wire [(9)-1:0] i_rtl_rstnn_seqeunce;
wire [(9)-1:0] i_rtl_rstpp_seqeunce;
wire i_rtl_rstnn_user;
wire i_rtl_rstpp_user;
wire [((1)*(1))-1:0] i_rtl_led_list;
wire i_rtl_i_xadc_wiz_0_clk;
wire i_rtl_i_xadc_wiz_0_rstnn;
wire i_rtl_i_system_ddr_clk_ref;
wire i_rtl_i_system_ddr_clk_sys;
wire i_rtl_i_system_ddr_rstnn_sys;
wire i_rtl_i_system_ddr_clk_dram_if;
wire i_rtl_i_system_ddr_rstnn_dram_if;
wire i_rtl_i_system_ddr_initialized;
wire i_rtl_i_pll0_external_rstnn;
wire i_rtl_i_pll0_clk_system;
wire i_rtl_i_pll0_clk_dram_sys;
wire i_rtl_i_pll0_clk_dram_ref;
wire i_rtl_i_system_sram_clk;
wire i_rtl_i_system_sram_rstnn;
wire [(1)-1:0] i_rtl_switch_slide_readymade_0_soe;
wire [(1)-1:0] i_rtl_switch_slide_readymade_0_soval;
wire [(1)-1:0] i_rtl_switch_slide_readymade_0_sival;
wire [(1)-1:0] i_rtl_gpio0_soe;
wire [(1)-1:0] i_rtl_gpio0_soval;
wire [(1)-1:0] i_rtl_gpio0_sival;
wire [(1)-1:0] i_rtl_gpio1_soe;
wire [(1)-1:0] i_rtl_gpio1_soval;
wire [(1)-1:0] i_rtl_gpio1_sival;
wire [(1)-1:0] i_rtl_gpio2_soe;
wire [(1)-1:0] i_rtl_gpio2_soval;
wire [(1)-1:0] i_rtl_gpio2_sival;
wire [(1)-1:0] i_rtl_gpio3_soe;
wire [(1)-1:0] i_rtl_gpio3_soval;
wire [(1)-1:0] i_rtl_gpio3_sival;
wire [(1)-1:0] i_rtl_gpio4_soe;
wire [(1)-1:0] i_rtl_gpio4_soval;
wire [(1)-1:0] i_rtl_gpio4_sival;
wire i_rtl_pjtag_rtck;
wire i_rtl_pjtag_rtrstnn;
wire i_rtl_pjtag_rtms;
wire i_rtl_pjtag_rtdi;
wire i_rtl_pjtag_rtdo;
wire i_rtl_printf_tx;
wire i_rtl_printf_rx;
wire i_rtl_i_xadc_wiz_0_sx4lawready;
wire i_rtl_i_xadc_wiz_0_sx4lawvalid;
wire [(32)-1:0] i_rtl_i_xadc_wiz_0_sx4lawaddr;
wire i_rtl_i_xadc_wiz_0_sx4lwready;
wire i_rtl_i_xadc_wiz_0_sx4lwvalid;
wire [(32)-1:0] i_rtl_i_xadc_wiz_0_sx4lwdata;
wire [(32/8)-1:0] i_rtl_i_xadc_wiz_0_sx4lwstrb;
wire i_rtl_i_xadc_wiz_0_sx4lbready;
wire i_rtl_i_xadc_wiz_0_sx4lbvalid;
wire [(2)-1:0] i_rtl_i_xadc_wiz_0_sx4lbresp;
wire i_rtl_i_xadc_wiz_0_sx4larready;
wire i_rtl_i_xadc_wiz_0_sx4larvalid;
wire [(32)-1:0] i_rtl_i_xadc_wiz_0_sx4laraddr;
wire i_rtl_i_xadc_wiz_0_sx4lrready;
wire i_rtl_i_xadc_wiz_0_sx4lrvalid;
wire [(32)-1:0] i_rtl_i_xadc_wiz_0_sx4lrdata;
wire [(2)-1:0] i_rtl_i_xadc_wiz_0_sx4lrresp;
wire i_rtl_i_system_ddr_sxawready;
wire i_rtl_i_system_ddr_sxawvalid;
wire [(32)-1:0] i_rtl_i_system_ddr_sxawaddr;
wire [(16)-1:0] i_rtl_i_system_ddr_sxawid;
wire [(8)-1:0] i_rtl_i_system_ddr_sxawlen;
wire [(3)-1:0] i_rtl_i_system_ddr_sxawsize;
wire [(2)-1:0] i_rtl_i_system_ddr_sxawburst;
wire i_rtl_i_system_ddr_sxwready;
wire i_rtl_i_system_ddr_sxwvalid;
wire [(16)-1:0] i_rtl_i_system_ddr_sxwid;
wire [(32)-1:0] i_rtl_i_system_ddr_sxwdata;
wire [(32/8)-1:0] i_rtl_i_system_ddr_sxwstrb;
wire i_rtl_i_system_ddr_sxwlast;
wire i_rtl_i_system_ddr_sxbready;
wire i_rtl_i_system_ddr_sxbvalid;
wire [(16)-1:0] i_rtl_i_system_ddr_sxbid;
wire [(2)-1:0] i_rtl_i_system_ddr_sxbresp;
wire i_rtl_i_system_ddr_sxarready;
wire i_rtl_i_system_ddr_sxarvalid;
wire [(32)-1:0] i_rtl_i_system_ddr_sxaraddr;
wire [(16)-1:0] i_rtl_i_system_ddr_sxarid;
wire [(8)-1:0] i_rtl_i_system_ddr_sxarlen;
wire [(3)-1:0] i_rtl_i_system_ddr_sxarsize;
wire [(2)-1:0] i_rtl_i_system_ddr_sxarburst;
wire i_rtl_i_system_ddr_sxrready;
wire i_rtl_i_system_ddr_sxrvalid;
wire [(16)-1:0] i_rtl_i_system_ddr_sxrid;
wire [(32)-1:0] i_rtl_i_system_ddr_sxrdata;
wire i_rtl_i_system_ddr_sxrlast;
wire [(2)-1:0] i_rtl_i_system_ddr_sxrresp;
wire i_rtl_i_system_sram_sxawready;
wire i_rtl_i_system_sram_sxawvalid;
wire [(32)-1:0] i_rtl_i_system_sram_sxawaddr;
wire [(`REQUIRED_BW_OF_SLAVE_TID)-1:0] i_rtl_i_system_sram_sxawid;
wire [(8)-1:0] i_rtl_i_system_sram_sxawlen;
wire [(3)-1:0] i_rtl_i_system_sram_sxawsize;
wire [(2)-1:0] i_rtl_i_system_sram_sxawburst;
wire i_rtl_i_system_sram_sxwready;
wire i_rtl_i_system_sram_sxwvalid;
wire [(`REQUIRED_BW_OF_SLAVE_TID)-1:0] i_rtl_i_system_sram_sxwid;
wire [(32)-1:0] i_rtl_i_system_sram_sxwdata;
wire [(32/8)-1:0] i_rtl_i_system_sram_sxwstrb;
wire i_rtl_i_system_sram_sxwlast;
wire i_rtl_i_system_sram_sxbready;
wire i_rtl_i_system_sram_sxbvalid;
wire [(`REQUIRED_BW_OF_SLAVE_TID)-1:0] i_rtl_i_system_sram_sxbid;
wire [(2)-1:0] i_rtl_i_system_sram_sxbresp;
wire i_rtl_i_system_sram_sxarready;
wire i_rtl_i_system_sram_sxarvalid;
wire [(32)-1:0] i_rtl_i_system_sram_sxaraddr;
wire [(`REQUIRED_BW_OF_SLAVE_TID)-1:0] i_rtl_i_system_sram_sxarid;
wire [(8)-1:0] i_rtl_i_system_sram_sxarlen;
wire [(3)-1:0] i_rtl_i_system_sram_sxarsize;
wire [(2)-1:0] i_rtl_i_system_sram_sxarburst;
wire i_rtl_i_system_sram_sxrready;
wire i_rtl_i_system_sram_sxrvalid;
wire [(`REQUIRED_BW_OF_SLAVE_TID)-1:0] i_rtl_i_system_sram_sxrid;
wire [(32)-1:0] i_rtl_i_system_sram_sxrdata;
wire i_rtl_i_system_sram_sxrlast;
wire [(2)-1:0] i_rtl_i_system_sram_sxrresp;
wire i_xadc_wiz_0_clk;
wire i_xadc_wiz_0_rstnn;
wire i_xadc_wiz_0_rx4lawready;
wire i_xadc_wiz_0_rx4lawvalid;
wire [(32)-1:0] i_xadc_wiz_0_rx4lawaddr;
wire i_xadc_wiz_0_rx4lwready;
wire i_xadc_wiz_0_rx4lwvalid;
wire [(32)-1:0] i_xadc_wiz_0_rx4lwdata;
wire [(32/8)-1:0] i_xadc_wiz_0_rx4lwstrb;
wire i_xadc_wiz_0_rx4lbready;
wire i_xadc_wiz_0_rx4lbvalid;
wire [(2)-1:0] i_xadc_wiz_0_rx4lbresp;
wire i_xadc_wiz_0_rx4larready;
wire i_xadc_wiz_0_rx4larvalid;
wire [(32)-1:0] i_xadc_wiz_0_rx4laraddr;
wire i_xadc_wiz_0_rx4lrready;
wire i_xadc_wiz_0_rx4lrvalid;
wire [(32)-1:0] i_xadc_wiz_0_rx4lrdata;
wire [(2)-1:0] i_xadc_wiz_0_rx4lrresp;
wire i_system_ddr_clk_ref;
wire i_system_ddr_clk_sys;
wire i_system_ddr_rstnn_sys;
wire i_system_ddr_clk_dram_if;
wire i_system_ddr_rstnn_dram_if;
wire i_system_ddr_initialized;
wire i_system_ddr_rxawready;
wire i_system_ddr_rxawvalid;
wire [(32)-1:0] i_system_ddr_rxawaddr;
wire [(16)-1:0] i_system_ddr_rxawid;
wire [(8)-1:0] i_system_ddr_rxawlen;
wire [(3)-1:0] i_system_ddr_rxawsize;
wire [(2)-1:0] i_system_ddr_rxawburst;
wire i_system_ddr_rxwready;
wire i_system_ddr_rxwvalid;
wire [(16)-1:0] i_system_ddr_rxwid;
wire [(32)-1:0] i_system_ddr_rxwdata;
wire [(32/8)-1:0] i_system_ddr_rxwstrb;
wire i_system_ddr_rxwlast;
wire i_system_ddr_rxbready;
wire i_system_ddr_rxbvalid;
wire [(16)-1:0] i_system_ddr_rxbid;
wire [(2)-1:0] i_system_ddr_rxbresp;
wire i_system_ddr_rxarready;
wire i_system_ddr_rxarvalid;
wire [(32)-1:0] i_system_ddr_rxaraddr;
wire [(16)-1:0] i_system_ddr_rxarid;
wire [(8)-1:0] i_system_ddr_rxarlen;
wire [(3)-1:0] i_system_ddr_rxarsize;
wire [(2)-1:0] i_system_ddr_rxarburst;
wire i_system_ddr_rxrready;
wire i_system_ddr_rxrvalid;
wire [(16)-1:0] i_system_ddr_rxrid;
wire [(32)-1:0] i_system_ddr_rxrdata;
wire i_system_ddr_rxrlast;
wire [(2)-1:0] i_system_ddr_rxrresp;
wire i_pll0_external_clk;
wire i_pll0_external_clk_pair;
wire i_pll0_external_rstnn;
wire i_pll0_clk_system;
wire i_pll0_clk_dram_sys;
wire i_pll0_clk_dram_ref;
wire i_system_sram_clk;
wire i_system_sram_rstnn;
wire i_system_sram_rxawready;
wire i_system_sram_rxawvalid;
wire [(32)-1:0] i_system_sram_rxawaddr;
wire [(`REQUIRED_BW_OF_SLAVE_TID)-1:0] i_system_sram_rxawid;
wire [(8)-1:0] i_system_sram_rxawlen;
wire [(3)-1:0] i_system_sram_rxawsize;
wire [(2)-1:0] i_system_sram_rxawburst;
wire i_system_sram_rxwready;
wire i_system_sram_rxwvalid;
wire [(`REQUIRED_BW_OF_SLAVE_TID)-1:0] i_system_sram_rxwid;
wire [(32)-1:0] i_system_sram_rxwdata;
wire [(32/8)-1:0] i_system_sram_rxwstrb;
wire i_system_sram_rxwlast;
wire i_system_sram_rxbready;
wire i_system_sram_rxbvalid;
wire [(`REQUIRED_BW_OF_SLAVE_TID)-1:0] i_system_sram_rxbid;
wire [(2)-1:0] i_system_sram_rxbresp;
wire i_system_sram_rxarready;
wire i_system_sram_rxarvalid;
wire [(32)-1:0] i_system_sram_rxaraddr;
wire [(`REQUIRED_BW_OF_SLAVE_TID)-1:0] i_system_sram_rxarid;
wire [(8)-1:0] i_system_sram_rxarlen;
wire [(3)-1:0] i_system_sram_rxarsize;
wire [(2)-1:0] i_system_sram_rxarburst;
wire i_system_sram_rxrready;
wire i_system_sram_rxrvalid;
wire [(`REQUIRED_BW_OF_SLAVE_TID)-1:0] i_system_sram_rxrid;
wire [(32)-1:0] i_system_sram_rxrdata;
wire i_system_sram_rxrlast;
wire [(2)-1:0] i_system_sram_rxrresp;
wire [((1)*(1))-1:0] tristate_buffer_for_switch_slide_readymade_0_roe_list;
wire [((1)*(1))-1:0] tristate_buffer_for_switch_slide_readymade_0_roval_list;
wire [((1)*(1))-1:0] tristate_buffer_for_switch_slide_readymade_0_rival_list;
wire [((1)*(1))-1:0] tristate_buffer_for_gpio0_roe_list;
wire [((1)*(1))-1:0] tristate_buffer_for_gpio0_roval_list;
wire [((1)*(1))-1:0] tristate_buffer_for_gpio0_rival_list;
wire [((1)*(1))-1:0] tristate_buffer_for_gpio1_roe_list;
wire [((1)*(1))-1:0] tristate_buffer_for_gpio1_roval_list;
wire [((1)*(1))-1:0] tristate_buffer_for_gpio1_rival_list;
wire [((1)*(1))-1:0] tristate_buffer_for_gpio2_roe_list;
wire [((1)*(1))-1:0] tristate_buffer_for_gpio2_roval_list;
wire [((1)*(1))-1:0] tristate_buffer_for_gpio2_rival_list;
wire [((1)*(1))-1:0] tristate_buffer_for_gpio3_roe_list;
wire [((1)*(1))-1:0] tristate_buffer_for_gpio3_roval_list;
wire [((1)*(1))-1:0] tristate_buffer_for_gpio3_rival_list;
wire [((1)*(1))-1:0] tristate_buffer_for_gpio4_roe_list;
wire [((1)*(1))-1:0] tristate_buffer_for_gpio4_roval_list;
wire [((1)*(1))-1:0] tristate_buffer_for_gpio4_rival_list;

FSD_V1_RTL
i_rtl
(
	.clk_system(i_rtl_clk_system),
	.clk_dca_core(i_rtl_clk_dca_core),
	.clk_core(i_rtl_clk_core),
	.clk_system_external(i_rtl_clk_system_external),
	.clk_system_debug(i_rtl_clk_system_debug),
	.clk_local_access(i_rtl_clk_local_access),
	.clk_process_000(i_rtl_clk_process_000),
	.clk_process_001(i_rtl_clk_process_001),
	.clk_dram_if(i_rtl_clk_dram_if),
	.clk_dram_sys(i_rtl_clk_dram_sys),
	.clk_dram_ref(i_rtl_clk_dram_ref),
	.clk_noc(i_rtl_clk_noc),
	.gclk_system(i_rtl_gclk_system),
	.gclk_dca_core(i_rtl_gclk_dca_core),
	.gclk_core(i_rtl_gclk_core),
	.gclk_system_external(i_rtl_gclk_system_external),
	.gclk_system_debug(i_rtl_gclk_system_debug),
	.gclk_local_access(i_rtl_gclk_local_access),
	.gclk_process_000(i_rtl_gclk_process_000),
	.gclk_process_001(i_rtl_gclk_process_001),
	.gclk_noc(i_rtl_gclk_noc),
	.tick_1us(i_rtl_tick_1us),
	.tick_62d5ms(i_rtl_tick_62d5ms),
	.tick_gpio(i_rtl_tick_gpio),
	.spi_common_sclk(i_rtl_spi_common_sclk),
	.spi_common_sdq0(i_rtl_spi_common_sdq0),
	.external_rstnn(i_rtl_external_rstnn),
	.global_rstnn(i_rtl_global_rstnn),
	.global_rstpp(i_rtl_global_rstpp),
	.rstnn_seqeunce(i_rtl_rstnn_seqeunce),
	.rstpp_seqeunce(i_rtl_rstpp_seqeunce),
	.rstnn_user(i_rtl_rstnn_user),
	.rstpp_user(i_rtl_rstpp_user),
	.led_list(i_rtl_led_list),
	.i_xadc_wiz_0_clk(i_rtl_i_xadc_wiz_0_clk),
	.i_xadc_wiz_0_rstnn(i_rtl_i_xadc_wiz_0_rstnn),
	.i_system_ddr_clk_ref(i_rtl_i_system_ddr_clk_ref),
	.i_system_ddr_clk_sys(i_rtl_i_system_ddr_clk_sys),
	.i_system_ddr_rstnn_sys(i_rtl_i_system_ddr_rstnn_sys),
	.i_system_ddr_clk_dram_if(i_rtl_i_system_ddr_clk_dram_if),
	.i_system_ddr_rstnn_dram_if(i_rtl_i_system_ddr_rstnn_dram_if),
	.i_system_ddr_initialized(i_rtl_i_system_ddr_initialized),
	.i_pll0_external_rstnn(i_rtl_i_pll0_external_rstnn),
	.i_pll0_clk_system(i_rtl_i_pll0_clk_system),
	.i_pll0_clk_dram_sys(i_rtl_i_pll0_clk_dram_sys),
	.i_pll0_clk_dram_ref(i_rtl_i_pll0_clk_dram_ref),
	.i_system_sram_clk(i_rtl_i_system_sram_clk),
	.i_system_sram_rstnn(i_rtl_i_system_sram_rstnn),
	.switch_slide_readymade_0_soe(i_rtl_switch_slide_readymade_0_soe),
	.switch_slide_readymade_0_soval(i_rtl_switch_slide_readymade_0_soval),
	.switch_slide_readymade_0_sival(i_rtl_switch_slide_readymade_0_sival),
	.gpio0_soe(i_rtl_gpio0_soe),
	.gpio0_soval(i_rtl_gpio0_soval),
	.gpio0_sival(i_rtl_gpio0_sival),
	.gpio1_soe(i_rtl_gpio1_soe),
	.gpio1_soval(i_rtl_gpio1_soval),
	.gpio1_sival(i_rtl_gpio1_sival),
	.gpio2_soe(i_rtl_gpio2_soe),
	.gpio2_soval(i_rtl_gpio2_soval),
	.gpio2_sival(i_rtl_gpio2_sival),
	.gpio3_soe(i_rtl_gpio3_soe),
	.gpio3_soval(i_rtl_gpio3_soval),
	.gpio3_sival(i_rtl_gpio3_sival),
	.gpio4_soe(i_rtl_gpio4_soe),
	.gpio4_soval(i_rtl_gpio4_soval),
	.gpio4_sival(i_rtl_gpio4_sival),
	.pjtag_rtck(i_rtl_pjtag_rtck),
	.pjtag_rtrstnn(i_rtl_pjtag_rtrstnn),
	.pjtag_rtms(i_rtl_pjtag_rtms),
	.pjtag_rtdi(i_rtl_pjtag_rtdi),
	.pjtag_rtdo(i_rtl_pjtag_rtdo),
	.printf_tx(i_rtl_printf_tx),
	.printf_rx(i_rtl_printf_rx),
	.i_xadc_wiz_0_sx4lawready(i_rtl_i_xadc_wiz_0_sx4lawready),
	.i_xadc_wiz_0_sx4lawvalid(i_rtl_i_xadc_wiz_0_sx4lawvalid),
	.i_xadc_wiz_0_sx4lawaddr(i_rtl_i_xadc_wiz_0_sx4lawaddr),
	.i_xadc_wiz_0_sx4lwready(i_rtl_i_xadc_wiz_0_sx4lwready),
	.i_xadc_wiz_0_sx4lwvalid(i_rtl_i_xadc_wiz_0_sx4lwvalid),
	.i_xadc_wiz_0_sx4lwdata(i_rtl_i_xadc_wiz_0_sx4lwdata),
	.i_xadc_wiz_0_sx4lwstrb(i_rtl_i_xadc_wiz_0_sx4lwstrb),
	.i_xadc_wiz_0_sx4lbready(i_rtl_i_xadc_wiz_0_sx4lbready),
	.i_xadc_wiz_0_sx4lbvalid(i_rtl_i_xadc_wiz_0_sx4lbvalid),
	.i_xadc_wiz_0_sx4lbresp(i_rtl_i_xadc_wiz_0_sx4lbresp),
	.i_xadc_wiz_0_sx4larready(i_rtl_i_xadc_wiz_0_sx4larready),
	.i_xadc_wiz_0_sx4larvalid(i_rtl_i_xadc_wiz_0_sx4larvalid),
	.i_xadc_wiz_0_sx4laraddr(i_rtl_i_xadc_wiz_0_sx4laraddr),
	.i_xadc_wiz_0_sx4lrready(i_rtl_i_xadc_wiz_0_sx4lrready),
	.i_xadc_wiz_0_sx4lrvalid(i_rtl_i_xadc_wiz_0_sx4lrvalid),
	.i_xadc_wiz_0_sx4lrdata(i_rtl_i_xadc_wiz_0_sx4lrdata),
	.i_xadc_wiz_0_sx4lrresp(i_rtl_i_xadc_wiz_0_sx4lrresp),
	.i_system_ddr_sxawready(i_rtl_i_system_ddr_sxawready),
	.i_system_ddr_sxawvalid(i_rtl_i_system_ddr_sxawvalid),
	.i_system_ddr_sxawaddr(i_rtl_i_system_ddr_sxawaddr),
	.i_system_ddr_sxawid(i_rtl_i_system_ddr_sxawid),
	.i_system_ddr_sxawlen(i_rtl_i_system_ddr_sxawlen),
	.i_system_ddr_sxawsize(i_rtl_i_system_ddr_sxawsize),
	.i_system_ddr_sxawburst(i_rtl_i_system_ddr_sxawburst),
	.i_system_ddr_sxwready(i_rtl_i_system_ddr_sxwready),
	.i_system_ddr_sxwvalid(i_rtl_i_system_ddr_sxwvalid),
	.i_system_ddr_sxwid(i_rtl_i_system_ddr_sxwid),
	.i_system_ddr_sxwdata(i_rtl_i_system_ddr_sxwdata),
	.i_system_ddr_sxwstrb(i_rtl_i_system_ddr_sxwstrb),
	.i_system_ddr_sxwlast(i_rtl_i_system_ddr_sxwlast),
	.i_system_ddr_sxbready(i_rtl_i_system_ddr_sxbready),
	.i_system_ddr_sxbvalid(i_rtl_i_system_ddr_sxbvalid),
	.i_system_ddr_sxbid(i_rtl_i_system_ddr_sxbid),
	.i_system_ddr_sxbresp(i_rtl_i_system_ddr_sxbresp),
	.i_system_ddr_sxarready(i_rtl_i_system_ddr_sxarready),
	.i_system_ddr_sxarvalid(i_rtl_i_system_ddr_sxarvalid),
	.i_system_ddr_sxaraddr(i_rtl_i_system_ddr_sxaraddr),
	.i_system_ddr_sxarid(i_rtl_i_system_ddr_sxarid),
	.i_system_ddr_sxarlen(i_rtl_i_system_ddr_sxarlen),
	.i_system_ddr_sxarsize(i_rtl_i_system_ddr_sxarsize),
	.i_system_ddr_sxarburst(i_rtl_i_system_ddr_sxarburst),
	.i_system_ddr_sxrready(i_rtl_i_system_ddr_sxrready),
	.i_system_ddr_sxrvalid(i_rtl_i_system_ddr_sxrvalid),
	.i_system_ddr_sxrid(i_rtl_i_system_ddr_sxrid),
	.i_system_ddr_sxrdata(i_rtl_i_system_ddr_sxrdata),
	.i_system_ddr_sxrlast(i_rtl_i_system_ddr_sxrlast),
	.i_system_ddr_sxrresp(i_rtl_i_system_ddr_sxrresp),
	.i_system_sram_sxawready(i_rtl_i_system_sram_sxawready),
	.i_system_sram_sxawvalid(i_rtl_i_system_sram_sxawvalid),
	.i_system_sram_sxawaddr(i_rtl_i_system_sram_sxawaddr),
	.i_system_sram_sxawid(i_rtl_i_system_sram_sxawid),
	.i_system_sram_sxawlen(i_rtl_i_system_sram_sxawlen),
	.i_system_sram_sxawsize(i_rtl_i_system_sram_sxawsize),
	.i_system_sram_sxawburst(i_rtl_i_system_sram_sxawburst),
	.i_system_sram_sxwready(i_rtl_i_system_sram_sxwready),
	.i_system_sram_sxwvalid(i_rtl_i_system_sram_sxwvalid),
	.i_system_sram_sxwid(i_rtl_i_system_sram_sxwid),
	.i_system_sram_sxwdata(i_rtl_i_system_sram_sxwdata),
	.i_system_sram_sxwstrb(i_rtl_i_system_sram_sxwstrb),
	.i_system_sram_sxwlast(i_rtl_i_system_sram_sxwlast),
	.i_system_sram_sxbready(i_rtl_i_system_sram_sxbready),
	.i_system_sram_sxbvalid(i_rtl_i_system_sram_sxbvalid),
	.i_system_sram_sxbid(i_rtl_i_system_sram_sxbid),
	.i_system_sram_sxbresp(i_rtl_i_system_sram_sxbresp),
	.i_system_sram_sxarready(i_rtl_i_system_sram_sxarready),
	.i_system_sram_sxarvalid(i_rtl_i_system_sram_sxarvalid),
	.i_system_sram_sxaraddr(i_rtl_i_system_sram_sxaraddr),
	.i_system_sram_sxarid(i_rtl_i_system_sram_sxarid),
	.i_system_sram_sxarlen(i_rtl_i_system_sram_sxarlen),
	.i_system_sram_sxarsize(i_rtl_i_system_sram_sxarsize),
	.i_system_sram_sxarburst(i_rtl_i_system_sram_sxarburst),
	.i_system_sram_sxrready(i_rtl_i_system_sram_sxrready),
	.i_system_sram_sxrvalid(i_rtl_i_system_sram_sxrvalid),
	.i_system_sram_sxrid(i_rtl_i_system_sram_sxrid),
	.i_system_sram_sxrdata(i_rtl_i_system_sram_sxrdata),
	.i_system_sram_sxrlast(i_rtl_i_system_sram_sxrlast),
	.i_system_sram_sxrresp(i_rtl_i_system_sram_sxrresp)
);

FSD_V1_SLOW_DRAM_00
i_system_ddr
(
	.clk_ref(i_system_ddr_clk_ref),
	.clk_sys(i_system_ddr_clk_sys),
	.rstnn_sys(i_system_ddr_rstnn_sys),
	.clk_dram_if(i_system_ddr_clk_dram_if),
	.rstnn_dram_if(i_system_ddr_rstnn_dram_if),
	.initialized(i_system_ddr_initialized),
	.rxawready(i_system_ddr_rxawready),
	.rxawvalid(i_system_ddr_rxawvalid),
	.rxawaddr(i_system_ddr_rxawaddr),
	.rxawid(i_system_ddr_rxawid),
	.rxawlen(i_system_ddr_rxawlen),
	.rxawsize(i_system_ddr_rxawsize),
	.rxawburst(i_system_ddr_rxawburst),
	.rxwready(i_system_ddr_rxwready),
	.rxwvalid(i_system_ddr_rxwvalid),
	.rxwid(i_system_ddr_rxwid),
	.rxwdata(i_system_ddr_rxwdata),
	.rxwstrb(i_system_ddr_rxwstrb),
	.rxwlast(i_system_ddr_rxwlast),
	.rxbready(i_system_ddr_rxbready),
	.rxbvalid(i_system_ddr_rxbvalid),
	.rxbid(i_system_ddr_rxbid),
	.rxbresp(i_system_ddr_rxbresp),
	.rxarready(i_system_ddr_rxarready),
	.rxarvalid(i_system_ddr_rxarvalid),
	.rxaraddr(i_system_ddr_rxaraddr),
	.rxarid(i_system_ddr_rxarid),
	.rxarlen(i_system_ddr_rxarlen),
	.rxarsize(i_system_ddr_rxarsize),
	.rxarburst(i_system_ddr_rxarburst),
	.rxrready(i_system_ddr_rxrready),
	.rxrvalid(i_system_ddr_rxrvalid),
	.rxrid(i_system_ddr_rxrid),
	.rxrdata(i_system_ddr_rxrdata),
	.rxrlast(i_system_ddr_rxrlast),
	.rxrresp(i_system_ddr_rxrresp)
	`include "slow_dram_cell_port_mapping.vh"
);

FSD_V1_CLOCK_PLL_0_01
i_pll0
(
	.external_clk(i_pll0_external_clk),
	.external_clk_pair(i_pll0_external_clk_pair),
	.external_rstnn(i_pll0_external_rstnn),
	.clk_system(i_pll0_clk_system),
	.clk_dram_sys(i_pll0_clk_dram_sys),
	.clk_dram_ref(i_pll0_clk_dram_ref)
);

FSD_V1_SRAM_AXI_02
i_system_sram
(
	.clk(i_system_sram_clk),
	.rstnn(i_system_sram_rstnn),
	.rxawready(i_system_sram_rxawready),
	.rxawvalid(i_system_sram_rxawvalid),
	.rxawaddr(i_system_sram_rxawaddr),
	.rxawid(i_system_sram_rxawid),
	.rxawlen(i_system_sram_rxawlen),
	.rxawsize(i_system_sram_rxawsize),
	.rxawburst(i_system_sram_rxawburst),
	.rxwready(i_system_sram_rxwready),
	.rxwvalid(i_system_sram_rxwvalid),
	.rxwid(i_system_sram_rxwid),
	.rxwdata(i_system_sram_rxwdata),
	.rxwstrb(i_system_sram_rxwstrb),
	.rxwlast(i_system_sram_rxwlast),
	.rxbready(i_system_sram_rxbready),
	.rxbvalid(i_system_sram_rxbvalid),
	.rxbid(i_system_sram_rxbid),
	.rxbresp(i_system_sram_rxbresp),
	.rxarready(i_system_sram_rxarready),
	.rxarvalid(i_system_sram_rxarvalid),
	.rxaraddr(i_system_sram_rxaraddr),
	.rxarid(i_system_sram_rxarid),
	.rxarlen(i_system_sram_rxarlen),
	.rxarsize(i_system_sram_rxarsize),
	.rxarburst(i_system_sram_rxarburst),
	.rxrready(i_system_sram_rxrready),
	.rxrvalid(i_system_sram_rxrvalid),
	.rxrid(i_system_sram_rxrid),
	.rxrdata(i_system_sram_rxrdata),
	.rxrlast(i_system_sram_rxrlast),
	.rxrresp(i_system_sram_rxrresp)
);

TRISTATE_BUFFER_OE
#(
	.NUM_DATA(1),
	.BW_DATA(1)
)
tristate_buffer_for_switch_slide_readymade_0
(
	.inout_port_list(switch_slide_readymade_0),
	.roe_list(tristate_buffer_for_switch_slide_readymade_0_roe_list),
	.roval_list(tristate_buffer_for_switch_slide_readymade_0_roval_list),
	.rival_list(tristate_buffer_for_switch_slide_readymade_0_rival_list)
);

TRISTATE_BUFFER_OE
#(
	.NUM_DATA(1),
	.BW_DATA(1)
)
tristate_buffer_for_gpio0
(
	.inout_port_list(gpio0),
	.roe_list(tristate_buffer_for_gpio0_roe_list),
	.roval_list(tristate_buffer_for_gpio0_roval_list),
	.rival_list(tristate_buffer_for_gpio0_rival_list)
);

TRISTATE_BUFFER_OE
#(
	.NUM_DATA(1),
	.BW_DATA(1)
)
tristate_buffer_for_gpio1
(
	.inout_port_list(gpio1),
	.roe_list(tristate_buffer_for_gpio1_roe_list),
	.roval_list(tristate_buffer_for_gpio1_roval_list),
	.rival_list(tristate_buffer_for_gpio1_rival_list)
);

TRISTATE_BUFFER_OE
#(
	.NUM_DATA(1),
	.BW_DATA(1)
)
tristate_buffer_for_gpio2
(
	.inout_port_list(gpio2),
	.roe_list(tristate_buffer_for_gpio2_roe_list),
	.roval_list(tristate_buffer_for_gpio2_roval_list),
	.rival_list(tristate_buffer_for_gpio2_rival_list)
);

TRISTATE_BUFFER_OE
#(
	.NUM_DATA(1),
	.BW_DATA(1)
)
tristate_buffer_for_gpio3
(
	.inout_port_list(gpio3),
	.roe_list(tristate_buffer_for_gpio3_roe_list),
	.roval_list(tristate_buffer_for_gpio3_roval_list),
	.rival_list(tristate_buffer_for_gpio3_rival_list)
);

TRISTATE_BUFFER_OE
#(
	.NUM_DATA(1),
	.BW_DATA(1)
)
tristate_buffer_for_gpio4
(
	.inout_port_list(gpio4),
	.roe_list(tristate_buffer_for_gpio4_roe_list),
	.roval_list(tristate_buffer_for_gpio4_roval_list),
	.rival_list(tristate_buffer_for_gpio4_rival_list)
);

assign i_rtl_external_rstnn = external_rstnn;
assign i_xadc_wiz_0_clk = i_rtl_i_xadc_wiz_0_clk;
assign i_xadc_wiz_0_rstnn = i_rtl_i_xadc_wiz_0_rstnn;
assign i_system_ddr_clk_ref = i_rtl_i_system_ddr_clk_ref;
assign i_system_ddr_clk_sys = i_rtl_i_system_ddr_clk_sys;
assign i_system_ddr_rstnn_sys = i_rtl_i_system_ddr_rstnn_sys;
assign i_rtl_i_system_ddr_clk_dram_if = i_system_ddr_clk_dram_if;
assign i_system_ddr_rstnn_dram_if = i_rtl_i_system_ddr_rstnn_dram_if;
assign i_rtl_i_system_ddr_initialized = i_system_ddr_initialized;
assign i_pll0_external_clk = external_clk_0;
assign i_pll0_external_clk_pair = external_clk_0_pair;
assign i_pll0_external_rstnn = i_rtl_i_pll0_external_rstnn;
assign i_rtl_i_pll0_clk_system = i_pll0_clk_system;
assign i_rtl_i_pll0_clk_dram_sys = i_pll0_clk_dram_sys;
assign i_rtl_i_pll0_clk_dram_ref = i_pll0_clk_dram_ref;
assign i_system_sram_clk = i_rtl_i_system_sram_clk;
assign i_system_sram_rstnn = i_rtl_i_system_sram_rstnn;
assign clk_system = i_rtl_clk_system;
assign clk_dca_core = i_rtl_clk_dca_core;
assign clk_core = i_rtl_clk_core;
assign clk_system_external = i_rtl_clk_system_external;
assign clk_system_debug = i_rtl_clk_system_debug;
assign clk_local_access = i_rtl_clk_local_access;
assign clk_process_000 = i_rtl_clk_process_000;
assign clk_process_001 = i_rtl_clk_process_001;
assign clk_dram_if = i_rtl_clk_dram_if;
assign clk_dram_sys = i_rtl_clk_dram_sys;
assign clk_dram_ref = i_rtl_clk_dram_ref;
assign clk_noc = i_rtl_clk_noc;
assign gclk_system = i_rtl_gclk_system;
assign gclk_dca_core = i_rtl_gclk_dca_core;
assign gclk_core = i_rtl_gclk_core;
assign gclk_system_external = i_rtl_gclk_system_external;
assign gclk_system_debug = i_rtl_gclk_system_debug;
assign gclk_local_access = i_rtl_gclk_local_access;
assign gclk_process_000 = i_rtl_gclk_process_000;
assign gclk_process_001 = i_rtl_gclk_process_001;
assign gclk_noc = i_rtl_gclk_noc;
assign tick_1us = i_rtl_tick_1us;
assign tick_62d5ms = i_rtl_tick_62d5ms;
assign tick_gpio = i_rtl_tick_gpio;
assign spi_common_sclk = i_rtl_spi_common_sclk;
assign spi_common_sdq0 = i_rtl_spi_common_sdq0;
assign global_rstnn = i_rtl_global_rstnn;
assign global_rstpp = i_rtl_global_rstpp;
assign rstnn_seqeunce = i_rtl_rstnn_seqeunce;
assign rstpp_seqeunce = i_rtl_rstpp_seqeunce;
assign rstnn_user = i_rtl_rstnn_user;
assign rstpp_user = i_rtl_rstpp_user;
assign led_list[1*(0+1)-1 -:1] = i_rtl_led_list[1*(0+1)-1 -:1];
assign tristate_buffer_for_switch_slide_readymade_0_roe_list[1*(0+1)-1 -:1] = i_rtl_switch_slide_readymade_0_soe;
assign tristate_buffer_for_switch_slide_readymade_0_roval_list[1*(0+1)-1 -:1] = i_rtl_switch_slide_readymade_0_soval;
assign i_rtl_switch_slide_readymade_0_sival = tristate_buffer_for_switch_slide_readymade_0_rival_list[1*(0+1)-1 -:1];
assign tristate_buffer_for_gpio0_roe_list[1*(0+1)-1 -:1] = i_rtl_gpio0_soe;
assign tristate_buffer_for_gpio0_roval_list[1*(0+1)-1 -:1] = i_rtl_gpio0_soval;
assign i_rtl_gpio0_sival = tristate_buffer_for_gpio0_rival_list[1*(0+1)-1 -:1];
assign tristate_buffer_for_gpio1_roe_list[1*(0+1)-1 -:1] = i_rtl_gpio1_soe;
assign tristate_buffer_for_gpio1_roval_list[1*(0+1)-1 -:1] = i_rtl_gpio1_soval;
assign i_rtl_gpio1_sival = tristate_buffer_for_gpio1_rival_list[1*(0+1)-1 -:1];
assign tristate_buffer_for_gpio2_roe_list[1*(0+1)-1 -:1] = i_rtl_gpio2_soe;
assign tristate_buffer_for_gpio2_roval_list[1*(0+1)-1 -:1] = i_rtl_gpio2_soval;
assign i_rtl_gpio2_sival = tristate_buffer_for_gpio2_rival_list[1*(0+1)-1 -:1];
assign tristate_buffer_for_gpio3_roe_list[1*(0+1)-1 -:1] = i_rtl_gpio3_soe;
assign tristate_buffer_for_gpio3_roval_list[1*(0+1)-1 -:1] = i_rtl_gpio3_soval;
assign i_rtl_gpio3_sival = tristate_buffer_for_gpio3_rival_list[1*(0+1)-1 -:1];
assign tristate_buffer_for_gpio4_roe_list[1*(0+1)-1 -:1] = i_rtl_gpio4_soe;
assign tristate_buffer_for_gpio4_roval_list[1*(0+1)-1 -:1] = i_rtl_gpio4_soval;
assign i_rtl_gpio4_sival = tristate_buffer_for_gpio4_rival_list[1*(0+1)-1 -:1];
assign i_rtl_pjtag_rtck = pjtag_rtck;
assign i_rtl_pjtag_rtrstnn = pjtag_rtrstnn;
assign i_rtl_pjtag_rtms = pjtag_rtms;
assign i_rtl_pjtag_rtdi = pjtag_rtdi;
assign pjtag_rtdo = i_rtl_pjtag_rtdo;
assign printf_tx = i_rtl_printf_tx;
assign i_rtl_printf_rx = printf_rx;
assign i_rtl_i_xadc_wiz_0_sx4lawready = i_xadc_wiz_0_rx4lawready;
assign i_xadc_wiz_0_rx4lawvalid = i_rtl_i_xadc_wiz_0_sx4lawvalid;
assign i_xadc_wiz_0_rx4lawaddr = i_rtl_i_xadc_wiz_0_sx4lawaddr;
assign i_rtl_i_xadc_wiz_0_sx4lwready = i_xadc_wiz_0_rx4lwready;
assign i_xadc_wiz_0_rx4lwvalid = i_rtl_i_xadc_wiz_0_sx4lwvalid;
assign i_xadc_wiz_0_rx4lwdata = i_rtl_i_xadc_wiz_0_sx4lwdata;
assign i_xadc_wiz_0_rx4lwstrb = i_rtl_i_xadc_wiz_0_sx4lwstrb;
assign i_xadc_wiz_0_rx4lbready = i_rtl_i_xadc_wiz_0_sx4lbready;
assign i_rtl_i_xadc_wiz_0_sx4lbvalid = i_xadc_wiz_0_rx4lbvalid;
assign i_rtl_i_xadc_wiz_0_sx4lbresp = i_xadc_wiz_0_rx4lbresp;
assign i_rtl_i_xadc_wiz_0_sx4larready = i_xadc_wiz_0_rx4larready;
assign i_xadc_wiz_0_rx4larvalid = i_rtl_i_xadc_wiz_0_sx4larvalid;
assign i_xadc_wiz_0_rx4laraddr = i_rtl_i_xadc_wiz_0_sx4laraddr;
assign i_xadc_wiz_0_rx4lrready = i_rtl_i_xadc_wiz_0_sx4lrready;
assign i_rtl_i_xadc_wiz_0_sx4lrvalid = i_xadc_wiz_0_rx4lrvalid;
assign i_rtl_i_xadc_wiz_0_sx4lrdata = i_xadc_wiz_0_rx4lrdata;
assign i_rtl_i_xadc_wiz_0_sx4lrresp = i_xadc_wiz_0_rx4lrresp;
assign i_rtl_i_system_ddr_sxawready = i_system_ddr_rxawready;
assign i_system_ddr_rxawvalid = i_rtl_i_system_ddr_sxawvalid;
assign i_system_ddr_rxawaddr = i_rtl_i_system_ddr_sxawaddr;
assign i_system_ddr_rxawid = i_rtl_i_system_ddr_sxawid;
assign i_system_ddr_rxawlen = i_rtl_i_system_ddr_sxawlen;
assign i_system_ddr_rxawsize = i_rtl_i_system_ddr_sxawsize;
assign i_system_ddr_rxawburst = i_rtl_i_system_ddr_sxawburst;
assign i_rtl_i_system_ddr_sxwready = i_system_ddr_rxwready;
assign i_system_ddr_rxwvalid = i_rtl_i_system_ddr_sxwvalid;
assign i_system_ddr_rxwid = i_rtl_i_system_ddr_sxwid;
assign i_system_ddr_rxwdata = i_rtl_i_system_ddr_sxwdata;
assign i_system_ddr_rxwstrb = i_rtl_i_system_ddr_sxwstrb;
assign i_system_ddr_rxwlast = i_rtl_i_system_ddr_sxwlast;
assign i_system_ddr_rxbready = i_rtl_i_system_ddr_sxbready;
assign i_rtl_i_system_ddr_sxbvalid = i_system_ddr_rxbvalid;
assign i_rtl_i_system_ddr_sxbid = i_system_ddr_rxbid;
assign i_rtl_i_system_ddr_sxbresp = i_system_ddr_rxbresp;
assign i_rtl_i_system_ddr_sxarready = i_system_ddr_rxarready;
assign i_system_ddr_rxarvalid = i_rtl_i_system_ddr_sxarvalid;
assign i_system_ddr_rxaraddr = i_rtl_i_system_ddr_sxaraddr;
assign i_system_ddr_rxarid = i_rtl_i_system_ddr_sxarid;
assign i_system_ddr_rxarlen = i_rtl_i_system_ddr_sxarlen;
assign i_system_ddr_rxarsize = i_rtl_i_system_ddr_sxarsize;
assign i_system_ddr_rxarburst = i_rtl_i_system_ddr_sxarburst;
assign i_system_ddr_rxrready = i_rtl_i_system_ddr_sxrready;
assign i_rtl_i_system_ddr_sxrvalid = i_system_ddr_rxrvalid;
assign i_rtl_i_system_ddr_sxrid = i_system_ddr_rxrid;
assign i_rtl_i_system_ddr_sxrdata = i_system_ddr_rxrdata;
assign i_rtl_i_system_ddr_sxrlast = i_system_ddr_rxrlast;
assign i_rtl_i_system_ddr_sxrresp = i_system_ddr_rxrresp;
assign i_rtl_i_system_sram_sxawready = i_system_sram_rxawready;
assign i_system_sram_rxawvalid = i_rtl_i_system_sram_sxawvalid;
assign i_system_sram_rxawaddr = i_rtl_i_system_sram_sxawaddr;
assign i_system_sram_rxawid = i_rtl_i_system_sram_sxawid;
assign i_system_sram_rxawlen = i_rtl_i_system_sram_sxawlen;
assign i_system_sram_rxawsize = i_rtl_i_system_sram_sxawsize;
assign i_system_sram_rxawburst = i_rtl_i_system_sram_sxawburst;
assign i_rtl_i_system_sram_sxwready = i_system_sram_rxwready;
assign i_system_sram_rxwvalid = i_rtl_i_system_sram_sxwvalid;
assign i_system_sram_rxwid = i_rtl_i_system_sram_sxwid;
assign i_system_sram_rxwdata = i_rtl_i_system_sram_sxwdata;
assign i_system_sram_rxwstrb = i_rtl_i_system_sram_sxwstrb;
assign i_system_sram_rxwlast = i_rtl_i_system_sram_sxwlast;
assign i_system_sram_rxbready = i_rtl_i_system_sram_sxbready;
assign i_rtl_i_system_sram_sxbvalid = i_system_sram_rxbvalid;
assign i_rtl_i_system_sram_sxbid = i_system_sram_rxbid;
assign i_rtl_i_system_sram_sxbresp = i_system_sram_rxbresp;
assign i_rtl_i_system_sram_sxarready = i_system_sram_rxarready;
assign i_system_sram_rxarvalid = i_rtl_i_system_sram_sxarvalid;
assign i_system_sram_rxaraddr = i_rtl_i_system_sram_sxaraddr;
assign i_system_sram_rxarid = i_rtl_i_system_sram_sxarid;
assign i_system_sram_rxarlen = i_rtl_i_system_sram_sxarlen;
assign i_system_sram_rxarsize = i_rtl_i_system_sram_sxarsize;
assign i_system_sram_rxarburst = i_rtl_i_system_sram_sxarburst;
assign i_system_sram_rxrready = i_rtl_i_system_sram_sxrready;
assign i_rtl_i_system_sram_sxrvalid = i_system_sram_rxrvalid;
assign i_rtl_i_system_sram_sxrid = i_system_sram_rxrid;
assign i_rtl_i_system_sram_sxrdata = i_system_sram_rxrdata;
assign i_rtl_i_system_sram_sxrlast = i_system_sram_rxrlast;
assign i_rtl_i_system_sram_sxrresp = i_system_sram_rxrresp;

`include "fsd_v1_user_region.vh"

`ifdef USE_ILA
`include "ila_description.vh"
`endif

endmodule