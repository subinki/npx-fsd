`ifndef __MUNOC_PROCESS_ID_H__
`define __MUNOC_PROCESS_ID_H__

`define PROCESS_ID_I_MNIM_I_MAIN_CORE_INST (0)
`define PROCESS_ID_I_MNIM_I_SUB_CORE_001_INST (1)
`define PROCESS_ID_I_MNIM_I_MAIN_CORE_DATA_C (0)
`define PROCESS_ID_I_MNIM_I_SUB_CORE_001_DATA_C (1)
`define PROCESS_ID_I_MNIM_I_MAIN_CORE_DATA_UC (0)
`define PROCESS_ID_I_MNIM_I_SUB_CORE_001_DATA_UC (1)

`endif