`ifndef __DCA_MATRIX_LSU_INST_H__
`define __DCA_MATRIX_LSU_INST_H__

`include "dca_matrix_info.vh"
`include "dca_module_memorymap_offset.vh"

`define BW_DCA_MATRIX_LSU_INST (`BW_DCA_MATRIX_LSU_INST_OPCODE+`BW_DCA_MATRIX_INFO_ALIGNED)

`define DCA_MATRIX_LSU_INST_OPCODE_READ 0

`endif
