// ****************************************************************************
// ****************************************************************************
// Copyright SoC Design Research Group, All rights reservxd.
// Electronics and Telecommunications Research Institute (ETRI)
// 
// THESE DOCUMENTS CONTAIN CONFIDENTIAL INFORMATION AND KNOWLEDGE
// WHICH IS THE PROPERTY OF ETRI. NO PART OF THIS PUBLICATION IS
// TO BE USED FOR ANY OTHER PURPOSE, AND THESE ARE NOT TO BE
// REPRODUCED, COPIED, DISCLOSED, TRANSMITTED, STORED IN A RETRIEVAL
// SYSTEM OR TRANSLATED INTO ANY OTHER HUMAN OR COMPUTER LANGUAGE,
// IN ANY FORM, BY ANY MEANS, IN WHOLE OR IN PART, WITHOUT THE
// COMPLETE PRIOR WRITTEN PERMISSION OF ETRI.
// ****************************************************************************
// 2025-11-05
// Kyuseung Han (han@etri.re.kr)
// ****************************************************************************
// ****************************************************************************

`include "ervp_global.vh"





module DCA_MODULE_00 
(
  dca_port_00,
  dca_port_02,
  dca_port_01,

  dca_port_03,
  dca_port_06,

  dca_port_12,
  dca_port_11,
  
  dca_port_10,
  dca_port_05,

  dca_port_08,
  dca_port_09,
  dca_port_04,
  dca_port_07
);





parameter DCA_GPARA_3 = 10;
parameter DCA_GPARA_2 = 10;
parameter DCA_GPARA_0 = 8;
parameter DCA_GPARA_1 = 8;

input wire dca_port_00;
input wire dca_port_02;
input wire dca_port_01;

input wire [DCA_GPARA_0-1:0] dca_port_03;
input wire [DCA_GPARA_1-1:0] dca_port_06;

input wire dca_port_12;
output wire dca_port_11;

output wire dca_port_10;
output wire dca_port_05;

output wire dca_port_08;
output wire dca_port_09;
output wire dca_port_04;
output wire dca_port_07;

localparam  DCA_LPARA_2 = 2;
localparam  DCA_LPARA_6 = 0;
localparam  DCA_LPARA_4 = 1;
localparam  DCA_LPARA_3 = 2;

reg [DCA_LPARA_2-1:0] dca_signal_04;
wire dca_signal_07;

localparam  DCA_LPARA_1 = DCA_GPARA_0;

reg [DCA_LPARA_1-1:0] dca_signal_01;
wire dca_signal_17;

wire dca_signal_14;
wire dca_signal_19;
wire [DCA_LPARA_1-1:0] dca_signal_15;
wire dca_signal_09;

localparam  DCA_LPARA_0 = DCA_GPARA_1 + 1;

reg [DCA_LPARA_0-1:0] dca_signal_20;
reg [DCA_LPARA_0-1:0] dca_signal_08;
wire dca_signal_05;
wire dca_signal_11;

wire dca_signal_06;
wire dca_signal_16;
wire [DCA_LPARA_0-1:0] dca_signal_03;
wire dca_signal_10;

localparam  DCA_LPARA_5 = `MAX(DCA_GPARA_2,DCA_GPARA_3);

wire dca_signal_00;
wire dca_signal_13;
wire [DCA_LPARA_5-1:0] dca_signal_02;

wire dca_signal_12;
wire dca_signal_18;

always@(posedge dca_port_00, negedge dca_port_02)
begin
  if(dca_port_02==0)
    dca_signal_04 <= DCA_LPARA_6;
  else if(dca_port_01)
  begin
    if(dca_port_11)
      dca_signal_04 <= DCA_LPARA_6;
    else if(dca_port_12)
      dca_signal_04 <= DCA_LPARA_3;
    else if(dca_signal_19)
      dca_signal_04 <= DCA_LPARA_4;
    else if(dca_signal_04==DCA_LPARA_4)
      dca_signal_04 <= DCA_LPARA_3;
  end
end

assign dca_signal_07 = (dca_signal_04==DCA_LPARA_3);

always@(posedge dca_port_00, negedge dca_port_02)
begin
  if(dca_port_02==0)
    dca_signal_01 <= 0;
  else if(dca_port_01)
  begin
    if(dca_port_12)
      dca_signal_01 <= dca_port_03;
    else if(dca_signal_19)
      dca_signal_01 <= (dca_signal_01>>1);
  end
end

assign dca_signal_17 = dca_signal_07 & dca_signal_01[0];

ERVP_COUNTER_WITH_ONEHOT_ENCODING
#(
  .COUNT_LENGTH(DCA_LPARA_1),
  .UP(1),
  .RESET_INDEX(0),
  .CIRCULAR(1)
)
i_dca_instance_1
(
  .clk(dca_port_00),
  .rstnn(dca_port_02),
  .enable(dca_port_01),
  .init(dca_signal_14),
  .count(dca_signal_19),
  .value(dca_signal_15),
  .is_first_count(),
  .is_last_count(dca_signal_09)
);

assign dca_signal_14 = dca_port_12;
assign dca_signal_19 = dca_signal_16 & dca_signal_10;

always@(posedge dca_port_00, negedge dca_port_02)
begin
  if(dca_port_02==0)
    dca_signal_20 <= 0;
  else if(dca_port_01)
  begin
    if(dca_port_12 || dca_signal_19)
      dca_signal_20 <= dca_port_06;
    else if(dca_signal_16)
      dca_signal_20 <= (dca_signal_20>>1);
  end
end

assign dca_signal_05 =  dca_signal_17 & dca_signal_20[0];

always@(posedge dca_port_00, negedge dca_port_02)
begin
  if(dca_port_02==0)
    dca_signal_08 <= 0;
  else if(dca_port_01)
  begin
    if(dca_port_12 || dca_signal_19)
      dca_signal_08 <= {dca_port_06,1'b 0};
    else if(dca_signal_16)
      dca_signal_08 <= (dca_signal_08>>1);
  end
end

assign dca_signal_11 = dca_signal_17 & dca_signal_08[0];

ERVP_COUNTER_WITH_ONEHOT_ENCODING
#(
  .COUNT_LENGTH(DCA_LPARA_0),
  .UP(1),
  .RESET_INDEX(0),
  .CIRCULAR(1)
)
i_dca_instance_2
(
  .clk(dca_port_00),
  .rstnn(dca_port_02),
  .enable(dca_port_01),
  .init(dca_signal_06),
  .count(dca_signal_16),
  .value(dca_signal_03),
  .is_first_count(),
  .is_last_count(dca_signal_10)
);

assign dca_signal_06 = dca_port_12 | dca_signal_19;
assign dca_signal_16 = dca_signal_07 & dca_signal_18;
assign dca_signal_12 = dca_signal_05 | dca_signal_11;
assign dca_signal_18 = dca_signal_12? dca_signal_02[DCA_LPARA_5-1] : 1;

ERVP_COUNTER_WITH_ONEHOT_ENCODING
#(
  .COUNT_LENGTH(DCA_LPARA_5),
  .UP(1),
  .RESET_INDEX(0),
  .CIRCULAR(1)
)
i_dca_instance_0
(
  .clk(dca_port_00),
  .rstnn(dca_port_02),
  .enable(dca_port_01),
  .init(dca_signal_00),
  .count(dca_signal_13),
  .value(dca_signal_02),
  .is_first_count(),
  .is_last_count()
);

assign dca_signal_00 = dca_port_12;
assign dca_signal_13 = dca_signal_12;

assign dca_port_10 = dca_signal_05 & dca_signal_02[0];
assign dca_port_05 = dca_signal_11 & dca_signal_02[0];

assign dca_port_11 = dca_signal_19 & dca_signal_09;

assign dca_port_08 = dca_signal_07 & dca_signal_10 & dca_signal_02[0];
assign dca_port_09 = dca_signal_07 & (~dca_signal_10) & dca_signal_02[0];
assign dca_port_04 = dca_signal_05 & dca_signal_02[DCA_GPARA_3-1];
assign dca_port_07 = dca_signal_11 & dca_signal_02[DCA_GPARA_2-1];

endmodule
